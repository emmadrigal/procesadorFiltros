module R_17_131071(output [16:0] o_reg);

assign o_reg=32'd131071;

endmodule 
