module DataMemory(input mem_WE,
						input mem_RE,
						input [31:0] Data,
						input [31:0] Dir,
						input clk,
						output [31:0] Data_out
						);

endmodule 