module R_4294967295(output [31:0] o_reg);

assign o_reg=32'd4294967295;

endmodule 