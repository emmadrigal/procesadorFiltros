module risk(input clk,
				input risk,
				input [3:0] OPCode,
				output ctrl,
				output atask
				);

endmodule 