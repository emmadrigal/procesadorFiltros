module adder(input [31:0]opA, input [31:0]opB, output[31:0] sum);

assign sum=opA+opB;

endmodule 