module Register(output [31:0] o_reg);

assign o_reg=32'd2;

endmodule 