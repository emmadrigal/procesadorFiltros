module R_16_65535(output [15:0] o_reg);

assign o_reg=32'd65535;

endmodule 