module Mem_Instructions( 
			input [31:0] i_dir,
			input clk,
			output [15:0] o_dir
			);

reg [15:0] mem_inst [0:255]; //[wordsize:0] a [0:arraysize]
reg [15:0] reg_o_dir;

reg initialized = 0;
reg done = 0;

always@(negedge clk) begin
	if(initialized == 0) begin
		mem_inst[0] <= 16'hb300;
		mem_inst[1] <= 16'hb200;
		mem_inst[2] <= 16'hb100;
		mem_inst[3] <= 16'h8b11;
		mem_inst[4] <= 16'he001;
		mem_inst[5] <= 16'hb30f;
		mem_inst[6] <= 16'hffff;
		mem_inst[7] <= 16'hb203;
		mem_inst[8] <= 16'hffff;
		mem_inst[9] <= 16'hffff;
		mem_inst[10] <= 16'hffff;
		mem_inst[11] <= 16'hffff;
		mem_inst[12] <= 16'hffff;
		mem_inst[13] <= 16'hffff;
		mem_inst[14] <= 16'hffff;
		mem_inst[15] <= 16'hffff;
		mem_inst[16] <= 16'hffff;
		mem_inst[17] <= 16'hffff;
		mem_inst[18] <= 16'hffff;
		mem_inst[19] <= 16'hffff;
		mem_inst[20] <= 16'hffff;
		mem_inst[21] <= 16'hffff;
		mem_inst[22] <= 16'hffff;
		mem_inst[23] <= 16'hffff;
		mem_inst[24] <= 16'hffff;
		mem_inst[25] <= 16'hffff;
		mem_inst[26] <= 16'hffff;
		mem_inst[27] <= 16'hffff;
		mem_inst[28] <= 16'hffff;
		mem_inst[29] <= 16'hffff;
		mem_inst[30] <= 16'hffff;
		mem_inst[31] <= 16'hffff;
		mem_inst[32] <= 16'hffff;
		mem_inst[33] <= 16'hffff;
		mem_inst[34] <= 16'hffff;
		mem_inst[35] <= 16'hffff;
		mem_inst[36] <= 16'hffff;
		mem_inst[37] <= 16'hffff;
		mem_inst[38] <= 16'hffff;
		mem_inst[39] <= 16'hffff;
		mem_inst[40] <= 16'hffff;
		mem_inst[41] <= 16'hffff;
		mem_inst[42] <= 16'hffff;
		mem_inst[43] <= 16'hffff;
		mem_inst[44] <= 16'hffff;
		mem_inst[45] <= 16'hffff;
		mem_inst[46] <= 16'hffff;
		mem_inst[47] <= 16'hffff;
		mem_inst[48] <= 16'hffff;
		mem_inst[49] <= 16'hffff;
		mem_inst[50] <= 16'hffff;
		mem_inst[51] <= 16'hffff;
		mem_inst[52] <= 16'hffff;
		mem_inst[53] <= 16'hffff;
		mem_inst[54] <= 16'hffff;
		mem_inst[55] <= 16'hffff;
		mem_inst[56] <= 16'hffff;
		mem_inst[57] <= 16'hffff;
		mem_inst[58] <= 16'hffff;
		mem_inst[59] <= 16'hffff;
		mem_inst[60] <= 16'hffff;
		mem_inst[61] <= 16'hffff;
		mem_inst[62] <= 16'hffff;
		mem_inst[63] <= 16'hffff;
		mem_inst[64] <= 16'hffff;
		mem_inst[65] <= 16'hffff;
		mem_inst[66] <= 16'hffff;
		mem_inst[67] <= 16'hffff;
		mem_inst[68] <= 16'hffff;
		mem_inst[69] <= 16'hffff;
		mem_inst[70] <= 16'hffff;
		mem_inst[71] <= 16'hffff;
		mem_inst[72] <= 16'hffff;
		mem_inst[73] <= 16'hffff;
		mem_inst[74] <= 16'hffff;
		mem_inst[75] <= 16'hffff;
		mem_inst[76] <= 16'hffff;
		mem_inst[77] <= 16'hffff;
		mem_inst[78] <= 16'hffff;
		mem_inst[79] <= 16'hffff;
		mem_inst[80] <= 16'hffff;
		mem_inst[81] <= 16'hffff;
		mem_inst[82] <= 16'hffff;
		mem_inst[83] <= 16'hffff;
		mem_inst[84] <= 16'hffff;
		mem_inst[85] <= 16'hffff;
		mem_inst[86] <= 16'hffff;
		mem_inst[87] <= 16'hffff;
		mem_inst[88] <= 16'hffff;
		mem_inst[89] <= 16'hffff;
		mem_inst[90] <= 16'hffff;
		mem_inst[91] <= 16'hffff;
		mem_inst[92] <= 16'hffff;
		mem_inst[93] <= 16'hffff;
		mem_inst[94] <= 16'hffff;
		mem_inst[95] <= 16'hffff;
		mem_inst[96] <= 16'hffff;
		mem_inst[97] <= 16'hffff;
		mem_inst[98] <= 16'hffff;
		mem_inst[99] <= 16'hffff;
		mem_inst[100] <= 16'hffff;
		mem_inst[101] <= 16'hffff;
		mem_inst[102] <= 16'hffff;
		mem_inst[103] <= 16'hffff;
		mem_inst[104] <= 16'hffff;
		mem_inst[105] <= 16'hffff;
		mem_inst[106] <= 16'hffff;
		mem_inst[107] <= 16'hffff;
		mem_inst[108] <= 16'hffff;
		mem_inst[109] <= 16'hffff;
		mem_inst[110] <= 16'hffff;
		mem_inst[111] <= 16'hffff;
		mem_inst[112] <= 16'hffff;
		mem_inst[113] <= 16'hffff;
		mem_inst[114] <= 16'hffff;
		mem_inst[115] <= 16'hffff;
		mem_inst[116] <= 16'hffff;
		mem_inst[117] <= 16'hffff;
		mem_inst[118] <= 16'hffff;
		mem_inst[119] <= 16'hffff;
		mem_inst[120] <= 16'hffff;
		mem_inst[121] <= 16'hffff;
		mem_inst[122] <= 16'hffff;
		mem_inst[123] <= 16'hffff;
		mem_inst[124] <= 16'hffff;
		mem_inst[125] <= 16'hffff;
		mem_inst[126] <= 16'hffff;
		mem_inst[127] <= 16'hffff;
		mem_inst[128] <= 16'hffff;
		mem_inst[129] <= 16'hffff;
		mem_inst[130] <= 16'hffff;
		mem_inst[131] <= 16'hffff;
		mem_inst[132] <= 16'hffff;
		mem_inst[133] <= 16'hffff;
		mem_inst[134] <= 16'hffff;
		mem_inst[135] <= 16'hffff;
		mem_inst[136] <= 16'hffff;
		mem_inst[137] <= 16'hffff;
		mem_inst[138] <= 16'hffff;
		mem_inst[139] <= 16'hffff;
		mem_inst[140] <= 16'hffff;
		mem_inst[141] <= 16'hffff;
		mem_inst[142] <= 16'hffff;
		mem_inst[143] <= 16'hffff;
		mem_inst[144] <= 16'hffff;
		mem_inst[145] <= 16'hffff;
		mem_inst[146] <= 16'hffff;
		mem_inst[147] <= 16'hffff;
		mem_inst[148] <= 16'hffff;
		mem_inst[149] <= 16'hffff;
		mem_inst[150] <= 16'hffff;
		mem_inst[151] <= 16'hffff;
		mem_inst[152] <= 16'hffff;
		mem_inst[153] <= 16'hffff;
		mem_inst[154] <= 16'hffff;
		mem_inst[155] <= 16'hffff;
		mem_inst[156] <= 16'hffff;
		mem_inst[157] <= 16'hffff;
		mem_inst[158] <= 16'hffff;
		mem_inst[159] <= 16'hffff;
		mem_inst[160] <= 16'hffff;
		mem_inst[161] <= 16'hffff;
		mem_inst[162] <= 16'hffff;
		mem_inst[163] <= 16'hffff;
		mem_inst[164] <= 16'hffff;
		mem_inst[165] <= 16'hffff;
		mem_inst[166] <= 16'hffff;
		mem_inst[167] <= 16'hffff;
		mem_inst[168] <= 16'hffff;
		mem_inst[169] <= 16'hffff;
		mem_inst[170] <= 16'hffff;
		mem_inst[171] <= 16'hffff;
		mem_inst[172] <= 16'hffff;
		mem_inst[173] <= 16'hffff;
		mem_inst[174] <= 16'hffff;
		mem_inst[175] <= 16'hffff;
		mem_inst[176] <= 16'hffff;
		mem_inst[177] <= 16'hffff;
		mem_inst[178] <= 16'hffff;
		mem_inst[179] <= 16'hffff;
		mem_inst[180] <= 16'hffff;
		mem_inst[181] <= 16'hffff;
		mem_inst[182] <= 16'hffff;
		mem_inst[183] <= 16'hffff;
		mem_inst[184] <= 16'hffff;
		mem_inst[185] <= 16'hffff;
		mem_inst[186] <= 16'hffff;
		mem_inst[187] <= 16'hffff;
		mem_inst[188] <= 16'hffff;
		mem_inst[189] <= 16'hffff;
		mem_inst[190] <= 16'hffff;
		mem_inst[191] <= 16'hffff;
		mem_inst[192] <= 16'hffff;
		mem_inst[193] <= 16'hffff;
		mem_inst[194] <= 16'hffff;
		mem_inst[195] <= 16'hffff;
		mem_inst[196] <= 16'hffff;
		mem_inst[197] <= 16'hffff;
		mem_inst[198] <= 16'hffff;
		mem_inst[199] <= 16'hffff;
		mem_inst[200] <= 16'hffff;
		mem_inst[201] <= 16'hffff;
		mem_inst[202] <= 16'hffff;
		mem_inst[203] <= 16'hffff;
		mem_inst[204] <= 16'hffff;
		mem_inst[205] <= 16'hffff;
		mem_inst[206] <= 16'hffff;
		mem_inst[207] <= 16'hffff;
		mem_inst[208] <= 16'hffff;
		mem_inst[209] <= 16'hffff;
		mem_inst[210] <= 16'hffff;
		mem_inst[211] <= 16'hffff;
		mem_inst[212] <= 16'hffff;
		mem_inst[213] <= 16'hffff;
		mem_inst[214] <= 16'hffff;
		mem_inst[215] <= 16'hffff;
		mem_inst[216] <= 16'hffff;
		mem_inst[217] <= 16'hffff;
		mem_inst[218] <= 16'hffff;
		mem_inst[219] <= 16'hffff;
		mem_inst[220] <= 16'hffff;
		mem_inst[221] <= 16'hffff;
		mem_inst[222] <= 16'hffff;
		mem_inst[223] <= 16'hffff;
		mem_inst[224] <= 16'hffff;
		mem_inst[225] <= 16'hffff;
		mem_inst[226] <= 16'hffff;
		mem_inst[227] <= 16'hffff;
		mem_inst[228] <= 16'hffff;
		mem_inst[229] <= 16'hffff;
		mem_inst[230] <= 16'hffff;
		mem_inst[231] <= 16'hffff;
		mem_inst[232] <= 16'hffff;
		mem_inst[233] <= 16'hffff;
		mem_inst[234] <= 16'hffff;
		mem_inst[235] <= 16'hffff;
		mem_inst[236] <= 16'hffff;
		mem_inst[237] <= 16'hffff;
		mem_inst[238] <= 16'hffff;
		mem_inst[239] <= 16'hffff;
		mem_inst[240] <= 16'hffff;
		mem_inst[241] <= 16'hffff;
		mem_inst[242] <= 16'hffff;
		mem_inst[243] <= 16'hffff;
		mem_inst[244] <= 16'hffff;
		mem_inst[245] <= 16'hffff;
		mem_inst[246] <= 16'hffff;
		mem_inst[247] <= 16'hffff;
		mem_inst[248] <= 16'hffff;
		mem_inst[249] <= 16'hffff;
		mem_inst[250] <= 16'hffff;
		mem_inst[251] <= 16'hffff;
		mem_inst[252] <= 16'hffff;
		mem_inst[253] <= 16'hffff;
		mem_inst[254] <= 16'hffff;
		mem_inst[255] <= 16'hffff;
		initialized <= 1;
	end
	
	if(i_dir == 255) begin
		done <= 1;
	end
	
	if(!done) begin
		reg_o_dir = mem_inst[i_dir];	
	end
end 


assign o_dir = reg_o_dir;


endmodule 