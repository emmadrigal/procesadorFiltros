module Register(output o_reg);

assign o_reg=32'd2;

endmodule 