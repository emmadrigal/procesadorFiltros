module ext(input [1:0] i,
				output [31:0] o
				);

endmodule 