module Truncate8(input [31:0] i,
					output [7:0] o
					);
					
assign o = i[7:0];

endmodule 