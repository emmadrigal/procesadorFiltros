module Register_Mem(input [3:0] DirA, 
						input [3:0] DirB, 
						input [3:0] Dir_WRA,  
						input [31:0]DI,	
						input clk,
						output [31:0]DatA, 
						output [31:0] DataB);

always@(posedge clk)begin

end

always@(negedge clk)begin

end

endmodule 