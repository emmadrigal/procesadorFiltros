module CMP_Combina(input ctrl,
						input [31:0] DatA,
						input [31:0] DatB,
						output risk
						);

endmodule 