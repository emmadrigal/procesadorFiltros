module R_1(output [31:0] o_reg);

assign o_reg=32'd1;

endmodule 