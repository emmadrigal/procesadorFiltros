module Regi(	input EN, 
			input [3:0] ia8,
			input [3:0] ib8,
			input [3:0] ic16,
			input [31:0] id32,
			input [31:0] ie32,
			input [31:0] if32,
			input [31:0] ig32,
			input [3:0] ih4,
			input [31:0] ij8,
			input clk,	
			
			output [3:0] oa8,
			output [3:0] ob8,
			output [3:0] oc16,
			output [31:0] od32,
			output [31:0] oe32,
			output [31:0] of32,
			output [31:0] og32,
			output [3:0] oh4,
			output [31:0] oj8
			);

endmodule 