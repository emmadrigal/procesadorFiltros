module ALU( input [3:0] code,
				input [31:0] X,
				input [31:0] Y,
				output [31:0] Z 
				);

endmodule 