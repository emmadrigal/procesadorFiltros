module R_32767(output [14:0] o_reg);

assign o_reg=32'd32767;

endmodule 