module Truncate4(input [31:0] i,
					output [3:0] o
);

assign o = i[3:0];

endmodule 