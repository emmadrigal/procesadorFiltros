module Ext8(input [7:0] i,
				output [31:0] o
				);

endmodule 